`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/17/2024 09:57:16 PM
// Design Name: 
// Module Name: tb_multiplier
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_multiplier();

    reg [31:0] a;
    reg [31:0] b;
    wire [31:0] p;
    
    // temp mantissa checking

    fp_multiplier uut (.num1(a), .num2(b), .final_product(p));
/*
    // mantissa checks
    initial begin
    
    #10 a = 32'd1;
    b = 32'd1;
    //100
    
    #10 a = 32'd3;
    b = 32'd3;
    //10000
    
    #10 a = 32'd7;
    b = 32'd7;
    //2730
    
    #10 a = 32'd15;
    b = 32'd15;
    //42435
    
    #10 a = 32'd31;
    b = 32'd31;
    
    
    #10 a = 32'd63;
    b = 32'd63;
    
    
    #10 a = 32'd127;
    b = 32'd127;
    
    
    #10 a = 32'd255;
    b = 32'd255;
    
    #10 a = 32'd511;
    b = 32'd511;
    
    #10 a = 32'd1023;
    b = 32'd1023;
    
    #10 a = 32'd2047;
    b = 32'd2047;
    
    #10 a = 32'd4095;
    b = 32'd4095;
    
    #10 a = 32'd8191;
    b = 32'd8191;
    
    
    
    end
    
    */
    initial begin
    
    // simple test of 1x1
    a = 32'b00111111100000000000000000000000; //1
    b = 32'b00111111100000000000000000000000; //1
    // expected result: same as above
    
    #30;
    // 2x2
    a = 32'b01000000000000000000000000000000;
    b = 32'b01000000000000000000000000000000;
    // expected result: 01000000100000000000000000000000
    
    #30;
    // 10x10
    a = 32'b01000001001000000000000000000000;
    b = 32'b01000001001000000000000000000000;
    
    
    #30;
    // 1.5x1.5
    a = 32'b00111111110000000000000000000000;
    b = 32'b00111111110000000000000000000000;
    
    #30;
    // 0.4x5
    a = 32'b00111110110011001100110011001101;
    b = 32'b01000000101000000000000000000000;
    
    #30;
    // 0x5
    a = 32'b00000000000000000000000000000000;
    b = 32'b01000000101000000000000000000000;
    
    #30;
    // 5x0
    a = 32'b01000000101000000000000000000000;
    b = 32'b00000000000000000000000000000000;
    
    #30;
    // 5xinf/NAN
    a = 32'b01000000101000000000000000000000;
    b = 32'b01111111100000000000000000000000;
    
    #30;
    // -inf/NANx5
    a = 32'b11111111100000000000000000000000;
    b = 32'b01000000101000000000000000000000;
    
    #30;
    // 12567x3490
    a = 32'b01000110010001000101110000000000;
    b = 32'b01000101010110100010000000000000;
    
    
    
    //0_100 0101 1_100 1000010100000000000
    //01000010100000000000000000000000
    
    
    // expected result: 01000010110010000000000000000000
    
    
    end
    

endmodule
